module not_gate(input logic a, output logic r);
    assign r = ~a;
endmodule
