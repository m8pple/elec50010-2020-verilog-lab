

module add_one(
    input logic[7:0] x,
    output logic[7:0] y
);

    assign y = x + 1;

endmodule